// alu_template.sv.j2
module alu_32bit (
    input  logic [31:0] A,
    input  logic [31:0] B,
    input  logic [2:0] opcode,
    output logic [31:0] result
);
    // Insert ALU logic here
endmodule